`default_nettype none

module instMemory(clk, reset, addr, inst);
  input wire clk, reset;
  input wire [31:0] addr;
  output logic [31:0] inst;

  (* ram_style = "block" *) 
  logic [31:0] mem [0:63];
  
  always_ff @(posedge clk) begin
    if(reset) begin
      mem[00] <= 32'b00001111110000000000010000010011;
      mem[01] <= 32'b00001101100000000000000100010011;
      mem[02] <= 32'b00000000000100010010101000100011;
      mem[03] <= 32'b00000000100000010010100000100011;
      mem[04] <= 32'b00000001110000010000010000010011;
      mem[05] <= 32'b00000000101000000000010100010011;
      mem[06] <= 32'b00000000110000000000000011101111;
      mem[07] <= 32'b00000000101000000010000000100011;
      mem[08] <= 32'b00000000000000000000000001101111;
      mem[09] <= 32'b00000000001001010010001010010011;
      mem[10] <= 32'b00000000000000101000011001100011;
      mem[11] <= 32'b00000000000100000000010100010011;
      mem[12] <= 32'b00000000000000001000000001100111;
      mem[13] <= 32'b11111110000000010000000100010011;
      mem[14] <= 32'b00000000000100010010101000100011;
      mem[15] <= 32'b00000000100000010010100000100011;
      mem[16] <= 32'b00000001110000010000010000010011;
      mem[17] <= 32'b00000000101001000010000000100011;
      mem[18] <= 32'b11111111111101010000010100010011;
      mem[19] <= 32'b11111101100111111111000011101111;
      mem[20] <= 32'b00000000101001000010001000100011;
      mem[21] <= 32'b00000000000001000010010100000011;
      mem[22] <= 32'b11111111111001010000010100010011;
      mem[23] <= 32'b11111100100111111111000011101111;
      mem[24] <= 32'b00000000010001000010010110000011;
      mem[25] <= 32'b00000000101101010000010100110011;
      mem[26] <= 32'b00000001010000010010000010000011;
      mem[27] <= 32'b00000001000000010010010000000011;
      mem[28] <= 32'b00000010000000010000000100010011;
      mem[29] <= 32'b00000000000000001000000001100111;
      for(int i=30; i<64; i=i+1) mem[i] <= 32'b0;
      inst <= 32'b00001111110000000000010000010011;
    end else begin
      inst <= mem[addr[7:2]];
    end
  end

endmodule

`default_nettype none